import uvm_pkg::*; // First import uvm_pkg then uvm_macros.svh
`include "uvm_macros.svh"
`include "jelly_bean_transaction.sv"
//import jelly_bean_pkg::*;
module top;
endmodule
